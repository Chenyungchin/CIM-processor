`timescale 1ns/10ps
`define CYCLE 10.0

module ReLU_tb;

// ================= clk generation =====================
reg clk = 1;
always #(`CYCLE/2) clk = ~clk;


// ================= dump waveform ======================
// vcd
initial begin
    $dumpfile("ReLU.vcd");
    $dumpvars(0, relu0);
end
// fsdb
// initial begin
//     $fsdbDumpfile("ReLu.fsdb");
//     $fsdbDumpvars(0, "+mda");
// end

// ================== time out ==========================
initial begin
    # (10000 * `CYCLE);
    $display("\n\033[1;31m=============================================");
	$display("           Simulation Time Out!      ");
	$display("=============================================\033[0m");
	$finish;
end

// ================= instantiate DUT ====================
parameter IN_PRECISION = 18;
parameter OUT_PRECISION = 4;
reg          rst_n = 1;
reg  [IN_PRECISION*64-1: 0]  relu_in;
wire [OUT_PRECISION*64-1: 0] relu_out;

ReLU #(
    .IN_PRECISION(IN_PRECISION),
    .OUT_PRECISION(OUT_PRECISION)
) relu0(
    .clk(clk),
    .rst_n(rst_n),
    .relu_in(relu_in),
    .relu_out(relu_out)
);


// ===== input pattern & result checking ===========
initial begin
    @(posedge clk) rst_n = 0;
    @(posedge clk) rst_n = 1;
    @(posedge clk) relu_in = 1152'b101010101010101010010101010101010101101010101010101010010101010101010101101010101010101010010101010101010101101010101010101010010101010101010101101010101010101010010101010101010101101010101010101010010101010101010101101010101010101010010101010101010101101010101010101010010101010101010101101010101010101010010101010101010101101010101010101010010101010101010101101010101010101010010101010101010101101010101010101010010101010101010101101010101010101010010101010101010101101010101010101010010101010101010101101010101010101010010101010101010101101010101010101010010101010101010101101010101010101010010101010101010101101010101010101010010101010101010101101010101010101010010101010101010101101010101010101010010101010101010101101010101010101010010101010101010101101010101010101010010101010101010101101010101010101010010101010101010101101010101010101010010101010101010101101010101010101010010101010101010101101010101010101010010101010101010101101010101010101010010101010101010101101010101010101010010101010101010101101010101010101010010101010101010101101010101010101010010101010101010101101010101010101010010101010101010101101010101010101010010101010101010101;
    @(posedge clk);
    @(posedge clk) relu_in = 1152'b010101010101010101101010101010101010010101010101010101101010101010101010010101010101010101101010101010101010010101010101010101101010101010101010010101010101010101101010101010101010010101010101010101101010101010101010010101010101010101101010101010101010010101010101010101101010101010101010010101010101010101101010101010101010010101010101010101101010101010101010010101010101010101101010101010101010010101010101010101101010101010101010010101010101010101101010101010101010010101010101010101101010101010101010010101010101010101101010101010101010010101010101010101101010101010101010010101010101010101101010101010101010010101010101010101101010101010101010010101010101010101101010101010101010010101010101010101101010101010101010010101010101010101101010101010101010010101010101010101101010101010101010010101010101010101101010101010101010010101010101010101101010101010101010010101010101010101101010101010101010010101010101010101101010101010101010010101010101010101101010101010101010010101010101010101101010101010101010010101010101010101101010101010101010010101010101010101101010101010101010010101010101010101101010101010101010010101010101010101101010101010101010;
    @(posedge clk);
    @(posedge clk);
    $finish;
end


endmodule