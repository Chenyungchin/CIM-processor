module Top(
    input    clk,
    input    rst_n,
    input    state,
    input    A,
    input    D,
    output   out_valid,
    output   Q
);



endmodule