// load data to mem
module LD(
    input    clk,
    input    rst_n,
    input [] act_in1_A,
    input [] act_in2_A,
    input [] act_in3_A,
    input [] weight_in_A,
    output [] act_in1,
    output [] act_in2,
    output [] act_in3,
    output [] weight_in
);

endmodule