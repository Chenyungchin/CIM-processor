module WB(
    input clk,
    input rst_n,
    input relu_out,
    input WB_A
);

endmodule